module token